module mycircuit( input logic [3:0]a, [2:0]s,
                  output logic seg_a, seg_b, seg_c, seg_d, seg_e, seg_f, seg_g, s1, s2, s3, s4, s5, s6, s7, s8  
);
assign seg_a = (~(a[3]) & ~(a[2]) & ~(a[1]) & a[0]) | (~(a[3]) & a[2] & ~(a[1]) & ~(a[0])) | (a[3] & a[2] & ~(a[1]) & a[0]) | (a[3] & ~(a[2]) & a[1] & a[0]);
assign seg_b = (~(a[3]) & a[2] & ~(a[1]) & a[0]) | (a[3] & a[2] & ~(a[1]) & ~(a[0])) | (a[2] & a[1] & ~(a[0])) | (a[3] & a[1] & a[0]);
assign seg_c = (a[3] & a[2] & ~(a[1]) & ~(a[0])) | (~(a[3]) & ~(a[2]) & a[1] & ~(a[0])) | (a[3] & a[2] & a[1]);
assign seg_d = (~(a[3]) & a[2] & ~(a[1]) & ~(a[0])) | (~(a[3]) & ~(a[2]) & ~(a[1]) & a[0]) | (a[2] & a[1] & a[0]) | (a[3] & ~(a[2]) & a[1] & ~(a[0]));  
assign seg_e = (~(a[3]) & a[2] & ~(a[1])) | (~(a[2]) & ~(a[1]) & a[0]) | (~(a[3]) & a[0]);
assign seg_f = (a[3] & a[2] & ~(a[1]) & a[0]) | (~(a[3]) & ~(a[2]) & a[0]) | (~(a[3]) & ~(a[2]) & a[1]) | (~(a[3]) & a[1] & a[0]);
assign seg_g = (~(a[3]) & ~(a[2]) & ~(a[1])) | (~(a[3]) & a[2] & a[1] & a[0]) | (a[3] & a[2] & ~(a[1]) & ~(a[0]));

assign s1 = (s[0] | s[1] | s[2]);
assign s2 = (~(s[0]) | s[1] | s[2]);
assign s3 = (s[0] | s[2] | ~(s[1]));
assign s4 = (~(s[0]) | s[2] | ~(s[1]));
assign s5 = (s[0] | ~(s[2]) | s[1]);
assign s6 = (~(s[0]) | ~(s[2]) | s[1]);
assign s7 = (s[0] | ~(s[2]) | ~(s[1]));
assign s8 = (~(s[0]) | ~(s[2]) | ~(s[1]));





endmodule